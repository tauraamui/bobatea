module bobatea

pub interface Contextable {}

struct Context {}

