module main

const shark_g = '🦈'
