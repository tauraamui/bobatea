module bobatea

import lib.draw

pub type Color = draw.Color
pub type Context = draw.Contextable
pub type Renderer = draw.Renderer
pub type Offset = draw.Offset
pub type ClipArea = draw.ClipArea
