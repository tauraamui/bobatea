module bobatea

import lib.draw

pub type Color = draw.Color
pub type Context = draw.Contextable
