// Copyright 2024 The Lilly Editor contributors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module draw

import lib.term.ui as tui

pub struct Event {
	tui.Event
}

pub struct Config {
pub:
	render_debug     bool
	default_fg_color ?Color
	default_bg_color ?Color
	user_data        voidptr
	frame_fn         fn (voidptr) @[required]
	update_fn        ?fn (voidptr) // Optional high-frequency update function
	event_fn         fn (Event, voidptr) @[required]

	capture_events       bool
	use_alternate_buffer bool = true
}

pub type Runner = fn () !

pub interface Drawer {
mut:
	set_stroke(s string)
	draw_text(x int, y int, text string)
	write(c string)
	draw_rect(x int, y int, width int, height int)
	draw_point(x int, y int)
	draw_line(x int, y int, x2 int, y2 int, do_apply_offsets bool)
}

pub interface Colorer {
mut:
	set_color(c Color)
	set_bg_color(c Color)
	set_default_fg_color(c Color)
	set_default_bg_color(c Color)
	get_default_fg_color() ?Color
	get_default_bg_color() ?Color
	reset_default_fg_color()
	reset_default_bg_color()
	reset_color()
	reset_bg_color()
}

pub interface Clipper {
mut:
	set_clip_area(c ClipArea)
	clear_clip_area()
}

pub interface WindowSizer {
	window_width() int
	window_height() int
}

pub interface Renderer {
	Drawer
	Colorer
	Clipper
	Offsetter
	WindowSizer
}

pub interface Contextable {
	Renderer
mut:
	render_debug() bool
	rate_limit_draws() bool

	set_cursor_position(x int, y int)
	set_cursor_to_block()
	set_cursor_to_underline()
	set_cursor_to_vertical_bar()
	show_cursor()
	hide_cursor()

	bold()
	set_style(s Style)
	clear_style()

	reset()

	//	run() !
	clear()
	flush()
	clear_prev_data()
}
